module test

endmodule
